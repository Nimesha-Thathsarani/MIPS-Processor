/*
    * CO224 - Computer Architecture
    * Lab 05 - Part 3
    * reg_file module
    * Version 1.0
*/

`include "cpu.v"

module Testbench;
    reg CLK, RESET;
    wire [31:0] PC;
    wire [31:0] INSTRUCTION;
    reg [7:0] instr_mem [0:1023];
    cpu mycpu(PC, INSTRUCTION, CLK, RESET);

    initial
    begin
        
        // METHOD 2: loading instr_mem content from instr_mem.mem file
        $readmemb("instr_mem.mem", instr_mem);
    end
    
    assign #2 INSTRUCTION ={instr_mem[PC+3] , instr_mem[PC+2] , instr_mem[PC+1],instr_mem[PC]};

    // always @ (PC)
    // begin
    //     # 2 // Latency for instruction register
    //     // Manually written opcodes

    //     case (PC)
    //     /*
    //         32'b0000_0000_0000_0000_0000_0000_0000_0000: INSTRUCTION = 32'b00000000_00000100_00000000_00000101; // loadi 4 0x05
            
    //         32'b0000_0000_0000_0000_0000_0000_0000_0100: INSTRUCTION = 32'b00000000_00000010_00000000_00001001; // loadi 2 0x09

    //         32'b0000_0000_0000_0000_0000_0000_0000_1000: INSTRUCTION = 32'b00000101_00000000_00000000_00000000; // add 6 4 2

    //         32'b0000_0000_0000_0000_0000_0000_0000_1100: INSTRUCTION = 32'b00000001_00000000_00000000_00000110; // mov 0 6
            
    //         32'b0000_0000_0000_0000_0000_0000_0001_0000: INSTRUCTION = 32'b00000000_00000001_00000000_00000001; // loadi 1 0x01
            
    //         32'b0000_0000_0000_0000_0000_0000_0001_0100: INSTRUCTION = 32'b00000010_00000010_00000010_00000001; // add 2 2 1

    //         32'b0000_0000_0000_0000_0000_0000_0001_1000: INSTRUCTION = 32'b00000110_00000000_00000000_00000000; // jmp 0
    //         */
            
    //         /*
    //         32'b0000_0000_0000_0000_0000_0000_0000_0000: INSTRUCTION = 32'b00000000_00000100_00000000_00000101; // loadi 4 0x05
            
    //         32'b0000_0000_0000_0000_0000_0000_0000_0100: INSTRUCTION = 32'b00000000_00000010_00000000_0000101; // loadi 2 0x09

    //         32'b0000_0000_0000_0000_0000_0000_0000_1000: INSTRUCTION = 32'b00000111_00000001_00000100_00000010; // add 6 4 2

    //         32'b0000_0000_0000_0000_0000_0000_0000_1100: INSTRUCTION = 32'b00000010_00000110_00000100_00000010; // mov 0 6
            
    //         32'b0000_0000_0000_0000_0000_0000_0001_0000: INSTRUCTION = 32'b00000000_00000110_00000000_00000011; // loadi 1 0x01
            
    //         32'b0000_0000_0000_0000_0000_0000_0001_0100: INSTRUCTION = 32'b00000001_00000000_00000000_00000110; // add 2 2 1

    //         32'b0000_0000_0000_0000_0000_0000_0001_1000: INSTRUCTION = 32'b00000110_00000001_00000000_00000000; // jmp 0

    //         32'b0000_0000_0000_0000_0000_0000_0001_1100: INSTRUCTION = 32'b00000000_00000001_00000000_00000001;

    //         32'b0000_0000_0000_0000_0000_0000_0010_0000: INSTRUCTION = 32'b00000010_00000010_00000010_00000000;

    //         */

    //         32'b0000_0000_0000_0000_0000_0000_0000_0000: INSTRUCTION = 32'b00000000_00000100_00000000_00001010; // loadi 4 0x05
            
    //         32'b0000_0000_0000_0000_0000_0000_0000_0100: INSTRUCTION = 32'b00000000_00000101_00000000_00000001; // loadi 2 0x09

    //         32'b0000_0000_0000_0000_0000_0000_0000_1000: INSTRUCTION = 32'b00000000_00000110_00000000_00000001; // add 6 4 2

    //         32'b0000_0000_0000_0000_0000_0000_0000_1100: INSTRUCTION = 32'b00000000_00000111_00000000_00001001; // mov 0 6
            
    //         32'b0000_0000_0000_0000_0000_0000_0001_0000: INSTRUCTION = 32'b00000011_00000100_00000100_00000101; // loadi 1 0x01
            
    //         32'b0000_0000_0000_0000_0000_0000_0001_0100: INSTRUCTION = 32'b00000111_00000001_00000100_00000110; // add 2 2 1

    //         32'b0000_0000_0000_0000_0000_0000_0001_1000: INSTRUCTION = 32'b00000110_11111101_00000000_00000000; // jmp 0

    //         32'b0000_0000_0000_0000_0000_0000_0001_1100: INSTRUCTION = 32'b00000010_00000001_00000100_00000111;

    //        // 32'b0000_0000_0000_0000_0000_0000_0010_0000: INSTRUCTION = 32'b00000010_00000010_00000010_00000000;
    //     endcase
    // end

    integer i;
    initial begin
        // generate files needed to plot the waveform using GTKWave
        $dumpfile("cpu_wavedata.vcd");
		$dumpvars(0, Testbench);
        
        for (i=0 ;i<8;i=i+1)
            $dumpvars(1,Testbench.mycpu.regfile.REGISTER[i]);
        
        
        RESET = 1'b0;
        CLK = 1'b0;
        
        // TODO: Reset the CPU (by giving a pulse to RESET signal) to start the program execution
        RESET = 1;
        #6
        RESET = 0;
        // finish simulation after some time
        #350
        $finish;
    end
        
    
    // clock signal generation
    always
        #4 CLK = ~CLK;
    
endmodule
module leftshift(
    input [31:0] data1,
    output [31:0] result
);

assign result=data1<<2;

endmodule

